////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//FSMpackageModule.sv - package module for output structre and enum value
//
//Author Prekshita Jain (prekjain@pdx.edu)
//date : 10/13/2018
//
//Description :
//______________________
// package module for output structre and enum value for states.
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
package FSMpackage;


typedef enum {READ1, IDLE} state;

typedef struct packed {
logic [7:0] data;
logic valid;
} out_st;

endpackage